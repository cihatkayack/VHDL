library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity frog_left_rom is
    Port (
        clk         : in  std_logic;
        address     : in  std_logic_vector(9 downto 0);
        color_data  : out std_logic_vector(11 downto 0)
    );
end frog_left_rom;

architecture Behavioral of frog_left_rom is
    type rom_type is array (0 to 783) of std_logic_vector(11 downto 0);
    signal rom : rom_type := (
        0 => "111111111111",
        1 => "111111111111",
        2 => "111111111111",
        3 => "111111111111",
        4 => "111111111111",
        5 => "000111110000",
        6 => "000111110000",
        7 => "111111111111",
        8 => "111111111111",
        9 => "111111111111",
        10 => "111111111111",
        11 => "111111111111",
        12 => "111111111111",
        13 => "111111111111",
        14 => "111111111111",
        15 => "111111111111",
        16 => "111111111111",
        17 => "111111111111",
        18 => "111111111111",
        19 => "111111111111",
        20 => "111111111111",
        21 => "000111110000",
        22 => "000111110000",
        23 => "111111111111",
        24 => "111111111111",
        25 => "111111111111",
        26 => "111111111111",
        27 => "111111111111",
        28 => "111111111111",
        29 => "111111111111",
        30 => "111111111111",
        31 => "111111111111",
        32 => "000111110000",
        33 => "000111110000",
        34 => "000111110000",
        35 => "000111110000",
        36 => "111111111111",
        37 => "111111111111",
        38 => "111111111111",
        39 => "111111111111",
        40 => "111111111111",
        41 => "111111111111",
        42 => "111111111111",
        43 => "111111111111",
        44 => "111111111111",
        45 => "111111111111",
        46 => "111111111111",
        47 => "111111111111",
        48 => "000111110000",
        49 => "000111110000",
        50 => "000111110000",
        51 => "000111110000",
        52 => "111111111111",
        53 => "111111111111",
        54 => "111111111111",
        55 => "111111111111",
        56 => "111111111111",
        57 => "111111111111",
        58 => "111111111111",
        59 => "111111111111",
        60 => "000111110000",
        61 => "000111110000",
        62 => "000111110000",
        63 => "000111110000",
        64 => "111111111111",
        65 => "111111111111",
        66 => "111111111111",
        67 => "111111111111",
        68 => "111111111111",
        69 => "111111111111",
        70 => "111111111111",
        71 => "111111111111",
        72 => "111111111111",
        73 => "111111111111",
        74 => "111111111111",
        75 => "111111111111",
        76 => "000111110000",
        77 => "000111110000",
        78 => "000111110000",
        79 => "000111110000",
        80 => "111111111111",
        81 => "111111111111",
        82 => "111111111111",
        83 => "111111111111",
        84 => "111111111111",
        85 => "000111110000",
        86 => "000111110000",
        87 => "000111110000",
        88 => "000111110000",
        89 => "000111110000",
        90 => "000111110000",
        91 => "000111110000",
        92 => "000111110000",
        93 => "000111110000",
        94 => "000111110000",
        95 => "111111111111",
        96 => "111111111111",
        97 => "111111111111",
        98 => "111111111111",
        99 => "111111111111",
        100 => "111111111111",
        101 => "000111110000",
        102 => "000111110000",
        103 => "000111110000",
        104 => "000111110000",
        105 => "000111110000",
        106 => "000111110000",
        107 => "000111110000",
        108 => "000111110000",
        109 => "000111110000",
        110 => "000111110000",
        111 => "111111111111",
        112 => "000111110000",
        113 => "000111110000",
        114 => "000111110000",
        115 => "000111110000",
        116 => "000111110000",
        117 => "000111110000",
        118 => "000111110000",
        119 => "000111110000",
        120 => "000111110000",
        121 => "000111110000",
        122 => "000111110000",
        123 => "000111110000",
        124 => "111111111111",
        125 => "111111111111",
        126 => "111111111111",
        127 => "111111111111",
        128 => "000111110000",
        129 => "000111110000",
        130 => "000111110000",
        131 => "000111110000",
        132 => "000111110000",
        133 => "000111110000",
        134 => "000111110000",
        135 => "000111110000",
        136 => "000111110000",
        137 => "000111110000",
        138 => "000111110000",
        139 => "000111110000",
        140 => "111111111111",
        141 => "000111110000",
        142 => "000111110000",
        143 => "000111110000",
        144 => "000111110000",
        145 => "000111110000",
        146 => "000111110000",
        147 => "000111110000",
        148 => "000111110000",
        149 => "000111110000",
        150 => "000111110000",
        151 => "000111110000",
        152 => "111111111111",
        153 => "111111111111",
        154 => "111111111111",
        155 => "111111111111",
        156 => "000111110000",
        157 => "000111110000",
        158 => "000111110000",
        159 => "000111110000",
        160 => "000111110000",
        161 => "000111110000",
        162 => "000111110000",
        163 => "000111110000",
        164 => "000111110000",
        165 => "000111110000",
        166 => "000111110000",
        167 => "111111111111",
        168 => "111111111111",
        169 => "111111111111",
        170 => "111111111111",
        171 => "111111111111",
        172 => "111111111111",
        173 => "111111111111",
        174 => "111111111111",
        175 => "111111111111",
        176 => "111111111111",
        177 => "000111110000",
        178 => "000111110000",
        179 => "000111110000",
        180 => "111111111111",
        181 => "111111111111",
        182 => "111111111111",
        183 => "111111111111",
        184 => "000111110000",
        185 => "000111110000",
        186 => "000111110000",
        187 => "111111111111",
        188 => "111111111111",
        189 => "111111111111",
        190 => "111111111111",
        191 => "111111111111",
        192 => "111111111111",
        193 => "111111111111",
        194 => "111111111111",
        195 => "111111111111",
        196 => "111111111111",
        197 => "111111111111",
        198 => "111111111111",
        199 => "111111111111",
        200 => "111111111111",
        201 => "111111111111",
        202 => "111111111111",
        203 => "111111111111",
        204 => "111111111111",
        205 => "000111110000",
        206 => "000111110000",
        207 => "000111110000",
        208 => "111111111111",
        209 => "111111111111",
        210 => "111111111111",
        211 => "111111111111",
        212 => "000111110000",
        213 => "000111110000",
        214 => "000111110000",
        215 => "111111111111",
        216 => "111111111111",
        217 => "111111111111",
        218 => "111111111111",
        219 => "111111111111",
        220 => "111111111111",
        221 => "111111111111",
        222 => "111111111111",
        223 => "111111111111",
        224 => "111111111111",
        225 => "111111111111",
        226 => "111111111111",
        227 => "111000001101",
        228 => "111000001101",
        229 => "000111110000",
        230 => "000111110000",
        231 => "111111110000",
        232 => "111111110000",
        233 => "111111110000",
        234 => "111111110000",
        235 => "111111110000",
        236 => "111111110000",
        237 => "111111110000",
        238 => "111111110000",
        239 => "111111110000",
        240 => "111111110000",
        241 => "111111110000",
        242 => "111111110000",
        243 => "111111110000",
        244 => "000111110000",
        245 => "111111111111",
        246 => "111111111111",
        247 => "111111111111",
        248 => "111111111111",
        249 => "111111111111",
        250 => "111111111111",
        251 => "111111111111",
        252 => "111111111111",
        253 => "111111111111",
        254 => "111000001101",
        255 => "111000001101",
        256 => "111000001101",
        257 => "000111110000",
        258 => "000111110000",
        259 => "111111110000",
        260 => "111111110000",
        261 => "000111110000",
        262 => "111111110000",
        263 => "111111110000",
        264 => "111111110000",
        265 => "111111110000",
        266 => "111111110000",
        267 => "111111110000",
        268 => "000111110000",
        269 => "111111110000",
        270 => "111111110000",
        271 => "111111110000",
        272 => "000111110000",
        273 => "000111110000",
        274 => "111111111111",
        275 => "111111111111",
        276 => "111111111111",
        277 => "111111111111",
        278 => "111111111111",
        279 => "111111111111",
        280 => "111111111111",
        281 => "111111111111",
        282 => "111000001101",
        283 => "111000001101",
        284 => "111000001101",
        285 => "000111110000",
        286 => "000111110000",
        287 => "111111110000",
        288 => "111111110000",
        289 => "000111110000",
        290 => "000111110000",
        291 => "111111110000",
        292 => "111111110000",
        293 => "111111110000",
        294 => "111111110000",
        295 => "000111110000",
        296 => "000111110000",
        297 => "111111110000",
        298 => "111111110000",
        299 => "111111110000",
        300 => "111111110000",
        301 => "000111110000",
        302 => "000111110000",
        303 => "111111111111",
        304 => "111111111111",
        305 => "111111111111",
        306 => "111111111111",
        307 => "111111111111",
        308 => "111111111111",
        309 => "111111110000",
        310 => "000111110000",
        311 => "000111110000",
        312 => "000111110000",
        313 => "000111110000",
        314 => "000111110000",
        315 => "111111110000",
        316 => "111111110000",
        317 => "111111110000",
        318 => "000111110000",
        319 => "000111110000",
        320 => "111111110000",
        321 => "111111110000",
        322 => "000111110000",
        323 => "111111110000",
        324 => "111111110000",
        325 => "111111110000",
        326 => "111111110000",
        327 => "111111110000",
        328 => "111111110000",
        329 => "111111110000",
        330 => "000111110000",
        331 => "000111110000",
        332 => "111111111111",
        333 => "111111111111",
        334 => "111111111111",
        335 => "111111111111",
        336 => "111111110000",
        337 => "111111110000",
        338 => "000111110000",
        339 => "000111110000",
        340 => "000111110000",
        341 => "000111110000",
        342 => "111111110000",
        343 => "111111110000",
        344 => "111111110000",
        345 => "111111110000",
        346 => "111111110000",
        347 => "000111110000",
        348 => "111111110000",
        349 => "111111110000",
        350 => "111111110000",
        351 => "111111110000",
        352 => "111111110000",
        353 => "111111110000",
        354 => "111111110000",
        355 => "111111110000",
        356 => "111111110000",
        357 => "111111110000",
        358 => "111111110000",
        359 => "111111110000",
        360 => "111111111111",
        361 => "111111111111",
        362 => "111111111111",
        363 => "111111111111",
        364 => "000111110000",
        365 => "111111110000",
        366 => "111111110000",
        367 => "111111110000",
        368 => "111111110000",
        369 => "111111110000",
        370 => "111111110000",
        371 => "111111110000",
        372 => "111111110000",
        373 => "111111110000",
        374 => "111111110000",
        375 => "111111110000",
        376 => "111111110000",
        377 => "111111110000",
        378 => "111111110000",
        379 => "111111110000",
        380 => "000111110000",
        381 => "000111110000",
        382 => "111111110000",
        383 => "111111110000",
        384 => "111111110000",
        385 => "111111110000",
        386 => "111111110000",
        387 => "111111110000",
        388 => "111111111111",
        389 => "111111111111",
        390 => "111111111111",
        391 => "111111111111",
        392 => "000111110000",
        393 => "111111110000",
        394 => "111111110000",
        395 => "111111110000",
        396 => "111111110000",
        397 => "111111110000",
        398 => "111111110000",
        399 => "111111110000",
        400 => "111111110000",
        401 => "111111110000",
        402 => "111111110000",
        403 => "111111110000",
        404 => "111111110000",
        405 => "111111110000",
        406 => "111111110000",
        407 => "000111110000",
        408 => "000111110000",
        409 => "000111110000",
        410 => "000111110000",
        411 => "111111110000",
        412 => "111111110000",
        413 => "111111110000",
        414 => "111111110000",
        415 => "111111110000",
        416 => "111111111111",
        417 => "111111111111",
        418 => "111111111111",
        419 => "111111111111",
        420 => "111111110000",
        421 => "111111110000",
        422 => "000111110000",
        423 => "000111110000",
        424 => "000111110000",
        425 => "000111110000",
        426 => "111111110000",
        427 => "111111110000",
        428 => "000111110000",
        429 => "111111110000",
        430 => "111111110000",
        431 => "111111110000",
        432 => "000111110000",
        433 => "000111110000",
        434 => "000111110000",
        435 => "000111110000",
        436 => "111111110000",
        437 => "111111110000",
        438 => "000111110000",
        439 => "000111110000",
        440 => "111111110000",
        441 => "111111110000",
        442 => "111111110000",
        443 => "111111110000",
        444 => "111111111111",
        445 => "111111111111",
        446 => "111111111111",
        447 => "111111111111",
        448 => "111111110000",
        449 => "111111110000",
        450 => "000111110000",
        451 => "000111110000",
        452 => "000111110000",
        453 => "000111110000",
        454 => "000111110000",
        455 => "111111110000",
        456 => "111111110000",
        457 => "000111110000",
        458 => "111111110000",
        459 => "111111110000",
        460 => "000111110000",
        461 => "000111110000",
        462 => "000111110000",
        463 => "000111110000",
        464 => "111111110000",
        465 => "111111110000",
        466 => "000111110000",
        467 => "000111110000",
        468 => "111111110000",
        469 => "111111110000",
        470 => "000111110000",
        471 => "000111110000",
        472 => "111111111111",
        473 => "111111111111",
        474 => "111111111111",
        475 => "111111111111",
        476 => "111111111111",
        477 => "111111111111",
        478 => "111000001101",
        479 => "111000001101",
        480 => "111000001101",
        481 => "000111110000",
        482 => "000111110000",
        483 => "111111110000",
        484 => "111111110000",
        485 => "000111110000",
        486 => "111111110000",
        487 => "111111110000",
        488 => "111111110000",
        489 => "111111110000",
        490 => "111111110000",
        491 => "000111110000",
        492 => "000111110000",
        493 => "000111110000",
        494 => "000111110000",
        495 => "111111110000",
        496 => "111111110000",
        497 => "000111110000",
        498 => "000111110000",
        499 => "111111111111",
        500 => "111111111111",
        501 => "111111111111",
        502 => "111111111111",
        503 => "111111111111",
        504 => "111111111111",
        505 => "111111111111",
        506 => "111000001101",
        507 => "111000001101",
        508 => "111000001101",
        509 => "000111110000",
        510 => "000111110000",
        511 => "111111110000",
        512 => "111111110000",
        513 => "111111110000",
        514 => "000111110000",
        515 => "111111110000",
        516 => "111111110000",
        517 => "111111110000",
        518 => "111111110000",
        519 => "111111110000",
        520 => "000111110000",
        521 => "000111110000",
        522 => "111111110000",
        523 => "111111110000",
        524 => "000111110000",
        525 => "000111110000",
        526 => "111111111111",
        527 => "111111111111",
        528 => "111111111111",
        529 => "111111111111",
        530 => "111111111111",
        531 => "111111111111",
        532 => "111111111111",
        533 => "111111111111",
        534 => "111111111111",
        535 => "111000001101",
        536 => "111000001101",
        537 => "000111110000",
        538 => "000111110000",
        539 => "111111110000",
        540 => "111111110000",
        541 => "111111110000",
        542 => "111111110000",
        543 => "111111110000",
        544 => "111111110000",
        545 => "111111110000",
        546 => "111111110000",
        547 => "111111110000",
        548 => "111111110000",
        549 => "111111110000",
        550 => "111111110000",
        551 => "000111110000",
        552 => "000111110000",
        553 => "111111111111",
        554 => "111111111111",
        555 => "111111111111",
        556 => "111111111111",
        557 => "111111111111",
        558 => "111111111111",
        559 => "111111111111",
        560 => "111111111111",
        561 => "111111111111",
        562 => "111111111111",
        563 => "111111111111",
        564 => "111111111111",
        565 => "111111111111",
        566 => "111111111111",
        567 => "111111111111",
        568 => "111111111111",
        569 => "000111110000",
        570 => "000111110000",
        571 => "000111110000",
        572 => "111111111111",
        573 => "111111111111",
        574 => "111111111111",
        575 => "111111111111",
        576 => "000111110000",
        577 => "000111110000",
        578 => "000111110000",
        579 => "111111111111",
        580 => "111111111111",
        581 => "111111111111",
        582 => "111111111111",
        583 => "111111111111",
        584 => "111111111111",
        585 => "111111111111",
        586 => "111111111111",
        587 => "111111111111",
        588 => "111111111111",
        589 => "111111111111",
        590 => "111111111111",
        591 => "111111111111",
        592 => "111111111111",
        593 => "111111111111",
        594 => "111111111111",
        595 => "111111111111",
        596 => "111111111111",
        597 => "000111110000",
        598 => "000111110000",
        599 => "000111110000",
        600 => "111111111111",
        601 => "111111111111",
        602 => "111111111111",
        603 => "111111111111",
        604 => "000111110000",
        605 => "000111110000",
        606 => "000111110000",
        607 => "111111111111",
        608 => "111111111111",
        609 => "111111111111",
        610 => "111111111111",
        611 => "111111111111",
        612 => "111111111111",
        613 => "111111111111",
        614 => "111111111111",
        615 => "111111111111",
        616 => "111111111111",
        617 => "000111110000",
        618 => "000111110000",
        619 => "000111110000",
        620 => "000111110000",
        621 => "000111110000",
        622 => "000111110000",
        623 => "000111110000",
        624 => "000111110000",
        625 => "000111110000",
        626 => "000111110000",
        627 => "000111110000",
        628 => "111111111111",
        629 => "111111111111",
        630 => "111111111111",
        631 => "111111111111",
        632 => "000111110000",
        633 => "000111110000",
        634 => "000111110000",
        635 => "000111110000",
        636 => "000111110000",
        637 => "000111110000",
        638 => "000111110000",
        639 => "000111110000",
        640 => "000111110000",
        641 => "000111110000",
        642 => "000111110000",
        643 => "111111111111",
        644 => "000111110000",
        645 => "000111110000",
        646 => "000111110000",
        647 => "000111110000",
        648 => "000111110000",
        649 => "000111110000",
        650 => "000111110000",
        651 => "000111110000",
        652 => "000111110000",
        653 => "000111110000",
        654 => "000111110000",
        655 => "000111110000",
        656 => "111111111111",
        657 => "111111111111",
        658 => "111111111111",
        659 => "111111111111",
        660 => "000111110000",
        661 => "000111110000",
        662 => "000111110000",
        663 => "000111110000",
        664 => "000111110000",
        665 => "000111110000",
        666 => "000111110000",
        667 => "000111110000",
        668 => "000111110000",
        669 => "000111110000",
        670 => "000111110000",
        671 => "000111110000",
        672 => "111111111111",
        673 => "000111110000",
        674 => "000111110000",
        675 => "000111110000",
        676 => "000111110000",
        677 => "000111110000",
        678 => "000111110000",
        679 => "000111110000",
        680 => "000111110000",
        681 => "000111110000",
        682 => "000111110000",
        683 => "111111111111",
        684 => "111111111111",
        685 => "111111111111",
        686 => "111111111111",
        687 => "111111111111",
        688 => "111111111111",
        689 => "000111110000",
        690 => "000111110000",
        691 => "000111110000",
        692 => "000111110000",
        693 => "000111110000",
        694 => "000111110000",
        695 => "000111110000",
        696 => "000111110000",
        697 => "000111110000",
        698 => "000111110000",
        699 => "111111111111",
        700 => "111111111111",
        701 => "111111111111",
        702 => "111111111111",
        703 => "111111111111",
        704 => "000111110000",
        705 => "000111110000",
        706 => "000111110000",
        707 => "000111110000",
        708 => "111111111111",
        709 => "111111111111",
        710 => "111111111111",
        711 => "111111111111",
        712 => "111111111111",
        713 => "111111111111",
        714 => "111111111111",
        715 => "111111111111",
        716 => "111111111111",
        717 => "111111111111",
        718 => "111111111111",
        719 => "111111111111",
        720 => "000111110000",
        721 => "000111110000",
        722 => "000111110000",
        723 => "000111110000",
        724 => "111111111111",
        725 => "111111111111",
        726 => "111111111111",
        727 => "111111111111",
        728 => "111111111111",
        729 => "111111111111",
        730 => "111111111111",
        731 => "111111111111",
        732 => "000111110000",
        733 => "000111110000",
        734 => "000111110000",
        735 => "000111110000",
        736 => "111111111111",
        737 => "111111111111",
        738 => "111111111111",
        739 => "111111111111",
        740 => "111111111111",
        741 => "111111111111",
        742 => "111111111111",
        743 => "111111111111",
        744 => "111111111111",
        745 => "111111111111",
        746 => "111111111111",
        747 => "111111111111",
        748 => "000111110000",
        749 => "000111110000",
        750 => "000111110000",
        751 => "000111110000",
        752 => "111111111111",
        753 => "111111111111",
        754 => "111111111111",
        755 => "111111111111",
        756 => "111111111111",
        757 => "111111111111",
        758 => "111111111111",
        759 => "111111111111",
        760 => "111111111111",
        761 => "000111110000",
        762 => "000111110000",
        763 => "111111111111",
        764 => "111111111111",
        765 => "111111111111",
        766 => "111111111111",
        767 => "111111111111",
        768 => "111111111111",
        769 => "111111111111",
        770 => "111111111111",
        771 => "111111111111",
        772 => "111111111111",
        773 => "111111111111",
        774 => "111111111111",
        775 => "111111111111",
        776 => "111111111111",
        777 => "000111110000",
        778 => "000111110000",
        779 => "111111111111",
        780 => "111111111111",
        781 => "111111111111",
        782 => "111111111111",
        783 => "111111111111"
    );
begin
    process(clk)
    begin
        if rising_edge(clk) then
            color_data <= rom(to_integer(unsigned(address)));
        end if;
    end process;
end Behavioral;
